grammar edu:umn:cs:melt:exts:ableC:regex:src ;

exports edu:umn:cs:melt:exts:ableC:regex:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:regex:src:concretesyntax ;